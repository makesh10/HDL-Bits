module top_module( input in, output out );
wire w;
    assign out=in;
endmodule
